.title KiCad schematic
.include "C:/AE/TLP183/B140HB.spice.txt"
.include "C:/AE/TLP183/ZR431.spice.txt"
.include "C:/AE/TLP183/c2012np02a102j060aa_p.mod"
.include "C:/AE/TLP183/c3216x5r1v106k160ab_p.mod"
.include "C:/AE/TLP183/TLP183.mod"
R4 /VOUT /VREF {RADJ}
R5 /VREF 0 {RREF}
XU3 /VZ /VCOMP C2012NP02A102J060AA_p
R3 /VCOMP /VREF {RCOMP}
I1 /VOUT 0 {ILOAD}
XU4 0 /VOUT C3216X5R1V106K160AB_p
V1 /VIN 0 {VSOURCE}
V2 /VC 0 {VSUPPLY}
R2 /VK /VZ {RZ}
R1 /VFB 0 {RE}
XU1 /VOUT /VK /VFB /VC TLP183
D1 /VIN /VOUT DI_B140HB
XU2 /VZ /VREF 0 ZR431
.end
